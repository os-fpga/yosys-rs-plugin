`include "./../SIM/SERDES_SIM/PLLTS16FFCFRACF.v"
`include "./../SIM/SERDES_SIM/PLLTS16FFCFRACF_library.v"
`include "./../SIM/SERDES_SIM/rs16.v"
`include "./../SIM/SERDES_SIM/rs_t16n20p90cpdlvt_ana.v"
`include "./../SIM/SERDES_SIM/phase_gen_4_8.v"
`include "./../SRC/GBX_SIM_MODEL_SRC/delay_line_tap64.sv"
`include "./../SRC/GBX_SIM_MODEL_SRC/phase_sel.sv"
`include "./../SRC/GBX_SIM_MODEL_SRC/gbox_bslip.sv"
`include "./../SRC/GBX_SIM_MODEL_SRC/gbox_cdr4.sv"
`include "./../SRC/GBX_SIM_MODEL_SRC/gbox_clk_gen.sv"
`include "./../SRC/GBX_SIM_MODEL_SRC/gbox_des.sv"
`include "./../SRC/GBX_SIM_MODEL_SRC/gbox_dly_adj.sv"
`include "./../SRC/GBX_SIM_MODEL_SRC/gbox_iobp_i.sv"
`include "./../SRC/GBX_SIM_MODEL_SRC/gbox_iobp_o.sv"
`include "./../SRC/GBX_SIM_MODEL_SRC/gbox_iobp_oe.sv"
`include "./../SRC/GBX_SIM_MODEL_SRC/gbox_rx.sv"
`include "./../SRC/GBX_SIM_MODEL_SRC/gbox_ser.sv"
`include "./../SRC/GBX_SIM_MODEL_SRC/gbox_top.sv"
`include "./../SRC/GBX_SIM_MODEL_SRC/gbox_tx.sv"
`include "./../SRC/GBX_SIM_MODEL_SRC/rs_sync_fifo_afe.sv"
`include "./../SRC/GBX_SIM_MODEL_SRC/rs_async_fifo_afe.v"
`include "./../SRC/GBX_SIM_MODEL_SRC/reset_sync.sv"
`include "./../SRC/GBX_SIM_MODEL_SRC/sync_flop.sv"


