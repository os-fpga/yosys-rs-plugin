`include "./../SRC/GBX/delay_line_tap64.sv"
`include "./../SRC/GBX/phase_sel.sv"
`include "./../SRC/GBX/gbox_bslip.sv"
`include "./../SRC/GBX/gbox_cdr4.sv"
`include "./../SRC/GBX/gbox_clk_gen.sv"
`include "./../SRC/GBX/gbox_des.sv"
`include "./../SRC/GBX/gbox_dly_adj.sv"
`include "./../SRC/GBX/gbox_iobp_i.sv"
`include "./../SRC/GBX/gbox_iobp_o.sv"
`include "./../SRC/GBX/gbox_iobp_oe.sv"
`include "./../SRC/GBX/gbox_rx.sv"
`include "./../SRC/GBX/gbox_ser.sv"
`include "./../SRC/GBX/gbox_top.sv"
`include "./../SRC/GBX/gbox_tx.sv"
`include "./../SRC/GBX/rs_sync_fifo_afe.sv"
`include "./../SRC/GBX/rs_async_fifo_afe.v"
`include "./../SRC/GBX/reset_sync.sv"
`include "./../SRC/GBX/sync_flop.sv"
